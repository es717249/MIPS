module Sim_Top_UartCtrl;




endmodule 