module TopMemory #(
	parameter DATA_WIDTH=32, 		//data length
	parameter ADDR_WIDTH=8			//bits to address the elements
)(

);