module TopMemory #(

)(

);